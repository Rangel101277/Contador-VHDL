library verilog;
use verilog.vl_types.all;
entity rangel_vlg_vec_tst is
end rangel_vlg_vec_tst;
